 `timescale 1ns / 1ps

module ALU(
    input [1:6] c,
    input [15:0] x,
    input [15:0] y,
    output [15:0] out,
    output zr,
    output ng
    );
    
// Your codes starts here

endmodule
